-- Package of utility functions for VHDL
-redacted:::




