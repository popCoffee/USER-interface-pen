-- package of procedures to support testing of VDP
-redacted::::



